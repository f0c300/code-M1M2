c<=b;
b<=a;
a<=a+b;
